*Title: Simple Verilog-A Resistor
.hdl resistor.va

.options post=1

X1 1 0 resistor r=1
VS 1 0 1

.dc VS 0 10 1

.end